interface intf;
  logic clk;
  logic rst;
  logic [2:0] count;
endinterface
