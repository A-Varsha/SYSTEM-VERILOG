// Code your testbench here
// or browse Examples
module associative_array_tb();
  associative_array dut();
  
  initial begin
    $dumpfile(associative_array.vcd);
    $dumpvars(0);
  end
endmodule
    
