# pass
#    monitor class signals      
# $time=16 rst=1 count =001
#        
# scb: not yet finished
# pass
#    monitor class signals      
# $time=36 rst=0 count =011
