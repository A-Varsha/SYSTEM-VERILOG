#       Generator        
# a=1 b=1 cin=0 sum=0 carry=0
#        
#        driver class signals         
# a=1 b=1 cin=0 sum=0 carry=0
#        
#       monitor class signals        
# a=1 b=1 cin=0 sum=0 carry=1
#        
# SCB: DUT=0/1 REF=0/1   PASS
#       monitor class signals        
# a=1 b=1 cin=0 sum=0 carry=1
#        
# SCB: DUT=0/1 REF=0/1   PASS
#       monitor class signals        
# a=1 b=1 cin=0 sum=0 carry=1
#        
# SCB: DUT=0/1 REF=0/1   PASS
#       monitor class signals        
# a=1 b=1 cin=0 sum=0 carry=1
#        
# SCB: DUT=0/1 REF=0/1   PASS
#       monitor class signals        
# a=1 b=1 cin=0 sum=0 carry=1
#        
# SCB: DUT=0/1 REF=0/1   PASS
#       Generator        
# a=1 b=1 cin=1 sum=0 carry=0
#        
#        driver class signals         
# a=1 b=1 cin=1 sum=0 carry=0
#        
#       Generator        
# a=0 b=1 cin=0 sum=0 carry=0
#        
#        driver class signals         
# a=0 b=1 cin=0 sum=0 carry=0
#        
#       Generator        
# a=1 b=0 cin=1 sum=0 carry=0
#        
#        driver class signals         
# a=1 b=0 cin=1 sum=0 carry=0
#        
#       Generator        
# a=1 b=1 cin=1 sum=0 carry=0
#        
#        driver class signals         
# a=1 b=1 cin=1 sum=0 carry=0
